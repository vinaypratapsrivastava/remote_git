module helloworld();
initial
begin
	$display (" this is first file Create");
	$display ("hello world");
	$display ("first modification");
end
endmodule
