module helloworld();
initial
begin
	$display (" this is first file Create");
	$display ("hello world");

end
endmodule
